//COMPILE: iverilog.exe -g2012 -o riscvsingle_p1.vcd -tvvp .\riscvsingle_p1.sv
//SIMULATE: vvp riscvsingle_p1


//------------------------------ TESTBENCH ------------------------//

module testbench();

  //Declara clock e reset com 1 bit
  logic        clk;
  logic        reset;

  //Declara WriteData e DataAdr com 32 bits e MemWrite com 1 bit
  logic [31:0] WriteData, DataAdr;
  logic        MemWrite;

  // instantiate device to be tested
  //Testa o modulo top clck e reset são inputs e o resto saida
  top dut(clk, reset, WriteData, DataAdr, MemWrite);
  
  // initialize test
  initial //Não repete
    begin
      reset <= 1; # 22; reset <= 0; //reset é 1 espera 22 tempos e reset fica 0
    end

  // generate clock to sequence tests
  always //Repete
    begin
      clk <= 1; # 5; clk <= 0; # 5; //Clock é 1 e depois de 5 tempos é 0
    end

  // check results
  always @(negedge clk) //Sempre no clock baixo
    begin
      if(MemWrite) //Só para ficar mais fácil de ver
        begin //Se MemWrite for 1 executa
          if(DataAdr === 100 && WriteData === 25) 
            begin //Se DataAdr for = 100 e WriteData = 25 //O === é para garantir sinais iguais //O & é para 1 bit
              $display("Simulation succeeded"); //Mostre isso
              $stop; //Pare
            end //Mesma coisa do begin
          else if (DataAdr !== 96) //Se DataAdr n for 96
            begin
              $display("Simulation failed");//Mostra isso
              $stop;//Para
            end
        end
    end
endmodule



//---------------------------------- COMEÇO DO CÓDIGO ----------------------------------------//


// ---- Instancia o processador, memória de dados e memória de instrução ---- //
//Cria o modulo do top
module top(input  logic        clk, reset, 
           output logic [31:0] WriteData, DataAdr, 
           output logic        MemWrite);//Clock e reset são inputs de 1 bit, WriteData e DataAdr são outputs de 32 bits, MemWrite é um output de 1 bit

  logic [31:0] PC, Instr, ReadData; //Cria o PC, Instr e ReadData com 32 bits
  
  // instantiate processor and memories
  //Cria rvsingle do tipo riscvsingle
  riscvsingle rvsingle(clk, reset, PC, Instr, MemWrite, DataAdr, 
                       WriteData, ReadData);//linha 78
  //cria imem do tipo imem
  imem imem(PC, Instr);
  //cria dmem do tipo dmem
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
endmodule



// --- Contém o controle e a lógica dos dados --- //
module riscvsingle(input  logic        clk, reset,//Clk e reset do top
                   output logic [31:0] PC,//Pc do top
                   input  logic [31:0] Instr,//Instr do top
                   output logic        MemWrite,//MemWrite do top
                   output logic [31:0] ALUResult, WriteData,//DataAdr e WriteData do top
                   input  logic [31:0] ReadData);//ReadData do top

  logic       ALUSrc, RegWrite, Jump, Zero;//Isso aí com 1 bit
  logic [1:0] ResultSrc, ImmSrc;//Isso aí com 2
  logic [2:0] ALUControl;//Isso aí com 3

  // Interpreta instrução e gera sinais de controle que ditam o comportamento. Lê os primeiros bits e decide a operação (add, sub, lw, etc) 
  //Usa o modulo controller
  controller c(Instr[6:0], Instr[14:12], Instr[30], Zero, 
               ResultSrc, MemWrite, PCSrc, 
               ALUSrc, RegWrite, Jump,
               ImmSrc, ALUControl);//linha 104
  
  // Manipulação dos dados durante execução. Unidades que fazem o cálculo real e acessam as memórias.
  datapath dp(clk, reset, ResultSrc, PCSrc,
              ALUSrc, RegWrite,
              ImmSrc, ALUControl,
              Zero, PC, Instr,
              ALUResult, WriteData, ReadData);
endmodule

module controller(input  logic [6:0] op,//Instr[6:0] do riscvsingle
                  input  logic [2:0] funct3,//Instr[14:12] do riscvsingle
                  input  logic       funct7b5,//Instr[30] do riscvsingle
                  input  logic       Zero,//Zero do riscvsingle
                  output logic [1:0] ResultSrc,//ResultSrc do riscvsingle
                  output logic       MemWrite,//MemWrite do riscvsingle
                  output logic       PCSrc, ALUSrc,//PCSrc e ALUSrc do riscvsingle
                  output logic       RegWrite, Jump,//RegWrite e jump do riscvsingle
                  output logic [1:0] ImmSrc,//ImmSrc do riscvsingle
                  output logic [2:0] ALUControl);//ALUControl do riscvsingle

  logic [1:0] ALUOp;
  logic       Branch;

  maindec md(op, ResultSrc, MemWrite, Branch,
             ALUSrc, RegWrite, Jump, ImmSrc, ALUOp);//126
  
  aludec  ad(op[5], funct3, funct7b5, ALUOp, ALUControl);

  assign PCSrc = Branch & Zero;
endmodule

module maindec(input  logic [6:0] op,
               output logic [1:0] ResultSrc,
               output logic       MemWrite,
               output logic       Branch, ALUSrc,
               output logic       RegWrite, Jump,
               output logic [1:0] ImmSrc,
               output logic [1:0] ALUOp);

  logic [10:0] controls;

  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp} = controls;

  always_comb
    case(op)
    // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
      7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type 
      7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
      default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // non-implemented instruction
    endcase
endmodule

module aludec(input  logic       opb5,
              input  logic [2:0] funct3,
              input  logic       funct7b5, 
              input  logic [1:0] ALUOp,
              output logic [2:0] ALUControl);

  logic  RtypeSub;
  assign RtypeSub = funct7b5 & opb5;  // TRUE for R-type subtract instruction

  always_comb
    case(ALUOp)
      2'b00:                ALUControl = 3'b000; // addition
      2'b01:                ALUControl = 3'b001; // subtraction
      default: case(funct3) // R-type or I-type ALU
                 3'b000:  if (RtypeSub) 
                            ALUControl = 3'b001; // sub
                          else          
                            ALUControl = 3'b000; // add, addi
                 3'b010:    ALUControl = 3'b101; // slt, slti
                 3'b110:    ALUControl = 3'b011; // or, ori
                 3'b111:    ALUControl = 3'b010; // and, andi
                 default:   ALUControl = 3'bxxx; // ???
               endcase
    endcase
endmodule

module datapath(input  logic        clk, reset,
                input  logic [1:0]  ResultSrc, 
                input  logic        PCSrc, ALUSrc,
                input  logic        RegWrite,
                input  logic [1:0]  ImmSrc,
                input  logic [2:0]  ALUControl,
                output logic        Zero,
                output logic [31:0] PC,
                input  logic [31:0] Instr,
                output logic [31:0] ALUResult, WriteData,
                input  logic [31:0] ReadData);

  logic [31:0] PCNext, PCPlus4, PCTarget;
  logic [31:0] ImmExt;
  logic [31:0] SrcA, SrcB;
  logic [31:0] Result;

  // next PC logic
  flopr #(32) pcreg(clk, reset, PCNext, PC); 
  adder       pcadd4(PC, 32'd4, PCPlus4);
  adder       pcaddbranch(PC, ImmExt, PCTarget);
  mux2 #(32)  pcmux(PCPlus4, PCTarget, PCSrc, PCNext);
 
  // register file logic
  regfile     rf(clk, RegWrite, Instr[19:15], Instr[24:20], 
                 Instr[11:7], Result, SrcA, WriteData);
  extend      ext(Instr[31:7], ImmSrc, ImmExt);

  // ALU logic
  mux2 #(32)  srcbmux(WriteData, ImmExt, ALUSrc, SrcB);
  alu         alu(SrcA, SrcB, ALUControl, ALUResult, Zero);
  mux3 #(32)  resultmux(ALUResult, ReadData, 32'b0, ResultSrc, Result);
endmodule


// --- Registradores de armazenamento temporário --- //
module regfile(input  logic        clk, 
               input  logic        we3, // a escrita ativa quando ele está alto
               input  logic [ 4:0] a1, a2, a3, // a1 e a2 servem para ler
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally (A1/RD1, A2/RD2)
  // write third port on rising edge of clock (A3/WD3/WE3)
  // register 0 hardwired to 0

  always_ff @(posedge clk)
    if (we3) rf[a3] <= wd3;	

  assign rd1 = (a1 != 0) ? rf[a1] : 0;
  assign rd2 = (a2 != 0) ? rf[a2] : 0;
endmodule

module adder(input  [31:0] a, b,
             output [31:0] y);

  assign y = a + b;
endmodule

module extend(input  logic [31:7] instr,
              input  logic [1:0]  immsrc,
              output logic [31:0] immext);
 
  always_comb
    case(immsrc) 
      2'b01:   immext = {{20{instr[31]}}, instr[31:25], instr[11:7]}; 
               // B-type (branches)
      2'b11:   immext = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0}; 
      default: immext = 32'bx; // undefined
    endcase             
endmodule

module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic             s, 
              output logic [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule

module mux3 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2,
              input  logic [1:0]       s, 
              output logic [WIDTH-1:0] y);

  assign y = s[1] ? d2 : (s[0] ? d1 : d0); 
endmodule

// --- Memória de instruções --- //
module imem(input  logic [31:0] a,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  initial
      $readmemh("riscvtest.txt",RAM);

  assign rd = RAM[a[31:2]]; // word aligned
endmodule

// --- Memória de dados --- //
module dmem(input  logic        clk, we,
            input  logic [31:0] a, wd,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  assign rd = RAM[a[31:2]]; // word aligned

  always_ff @(posedge clk)
    if (we) RAM[a[31:2]] <= wd;
endmodule




// --- Módulo da ALU --- //
module alu(input  logic [31:0] a, b,
           input  logic [2:0]  alucontrol,
           output logic [31:0] result,
           output logic        zero);

  logic [31:0] condinvb, sum;
  logic        v;              // overflow
  logic        isAddSub;       // true when is add or subtract operation

  
  //ALTERADO//
  
  assign zero = (result == 32'b0);// ESTAVA FORA DAS DECLARAÇÕES
  assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;// ESTAVA FORA DAS DECLARAÇÕES
  assign condinvb = alucontrol[0] ? ~b : b;
  assign sum = a + condinvb + alucontrol[0];
  assign isAddSub = ~alucontrol[2] & ~alucontrol[1] |
                    ~alucontrol[1] & alucontrol[0];

  always_comb
    case (alucontrol)
      3'b000:  result = sum;         // add
      3'b001:  result = sum;         // subtract
      3'b010:  result = a & b;       // and
      3'b011:  result = a | b;       // or
      3'b100:  result = a ^ b;       // xor
      3'b101:  result = sum[31] ^ v; // slt
      3'b110:  result = a << b[4:0]; // sll
      3'b111:  result = a >> b[4:0]; // srl
      default: result = 32'bx;
    endcase
  
endmodule

